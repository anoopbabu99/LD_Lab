module and16_gate(d,b,a);
input[15:0]a,b;
output[15:0]d;

and_gate and_gate_1[15:0](d,b,a);
endmodule 
