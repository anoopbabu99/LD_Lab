module stimulus;
wire s,c;
reg a,b;

halfadder halfadder_1(s,c,b,a);
initial 
begin

a=1'b0; b=1'b0;
#10 a=1'b0;b=1'b1; 
#10 a=1'b1;b=1'b0; 
#10 a=1'b1;b=1'b1;

end
endmodule
