module stimulus;
wire e;
reg a,b;


or_gate or_gate_1 (e,b,a);
initial
begin
a=1'b0; b=1'b0;
#10 a=1'b0;b=1'b1; 
#10 a=1'b1;b=1'b0; 
#10 a=1'b1;b=1'b1;
end
endmodule


