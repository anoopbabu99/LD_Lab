module stimulus;
wire a7,a6,a5,a4,a3,a2,a1,a0;
reg i,s2,s1,s0;

demux81_gate demux81_gate_1(i,s0,s1,s2,a7,a6,a5,a4,a3,a2,a1,a0);
initial
begin
i=1'b0; s2=1'b0; s1=1'b0; s0=1'b0;
#10 i=1'b0; s2=1'b0; s1=1'b0; s0=1'b1;
#10 i=1'b0; s2=1'b0; s1=1'b1; s0=1'b0;
#10 i=1'b0; s2=1'b0; s1=1'b1; s0=1'b1;
#10 i=1'b0; s2=1'b1; s1=1'b0; s0=1'b0;
#10 i=1'b0; s2=1'b1; s1=1'b0; s0=1'b1;
#10 i=1'b0; s2=1'b1; s1=1'b1; s0=1'b0;
#10 i=1'b0; s2=1'b1; s1=1'b1; s0=1'b1;
#10 i=1'b1; s2=1'b0; s1=1'b0; s0=1'b0;
#10 i=1'b1; s2=1'b0; s1=1'b0; s0=1'b1;
#10 i=1'b1; s2=1'b0; s1=1'b1; s0=1'b0;
#10 i=1'b1; s2=1'b0; s1=1'b1; s0=1'b1;
#10 i=1'b1; s2=1'b1; s1=1'b0; s0=1'b0;
#10 i=1'b1; s2=1'b1; s1=1'b0; s0=1'b1;
#10 i=1'b1; s2=1'b1; s1=1'b1; s0=1'b0;
#10 i=1'b1; s2=1'b1; s1=1'b1; s0=1'b1;

end
endmodule
